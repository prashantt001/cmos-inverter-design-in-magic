magic
tech scmos
timestamp 1660052862
<< polysilicon >>
rect 5 20 7 22
rect 5 -3 7 0
rect 3 -7 7 -3
rect 5 -10 7 -7
rect 5 -22 7 -20
<< ndiffusion >>
rect 4 -20 5 -10
rect 7 -20 8 -10
<< pdiffusion >>
rect 4 0 5 20
rect 7 0 8 20
<< metal1 >>
rect -4 28 16 29
rect -4 24 -3 28
rect 1 24 11 28
rect 15 24 16 28
rect -4 23 16 24
rect 0 20 4 23
rect 8 -10 12 0
rect 0 -23 4 -20
rect -4 -24 16 -23
rect -4 -28 -3 -24
rect 1 -28 11 -24
rect 15 -28 16 -24
rect -4 -29 16 -28
<< ntransistor >>
rect 5 -20 7 -10
<< ptransistor >>
rect 5 0 7 20
<< polycontact >>
rect -1 -7 3 -3
<< ndcontact >>
rect 0 -20 4 -10
rect 8 -20 12 -10
<< pdcontact >>
rect 0 0 4 20
rect 8 0 12 20
<< psubstratepcontact >>
rect -3 -28 1 -24
rect 11 -28 15 -24
<< nsubstratencontact >>
rect -3 24 1 28
rect 11 24 15 28
<< labels >>
rlabel metal1 3 25 3 25 5 vdd
rlabel metal1 3 -27 3 -27 1 gnd
rlabel metal1 10 -5 10 -5 1 Z
rlabel polycontact 1 -5 1 -5 3 A
<< end >>
